library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity char_rom is
    port(
        addr: in std_logic_vector(8 downto 0);
        data: out std_logic_vector(0 to 7)
    );
end char_rom;

architecture content of char_rom is
    type rom_type is array(0 to 335) of std_logic_vector(7 downto 0);
    constant FONT: rom_type :=
    (
        -- 0
        "00111000", -- ..###
        "01001100", -- .# .##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "01100100", -- .##..#
        "00111000", -- ..###
        "00000000", --
        -- 1 
        "00011000", -- ..##
        "00111000", -- .###
        "00011000", -- ..##
        "00011000", -- ..##
        "00011000", -- ..##
        "00011000", -- ..##
        "01111110", -- ######
        "00000000", --
        -- 2 
        "01111100", -- .#####
        "11000110", -- ##...##
        "00001110", -- ....###
        "00111100", -- ..####
        "01111000", -- .####
        "11100000", -- ###
        "11111110", -- #######
        "00000000", --
        -- 3 
        "01111110", -- .######
        "00001100", -- ....##
        "00011000", -- ...##
        "00111100", -- ..####
        "00000110", -- .....##
        "11000110", -- ##...##
        "01111100", -- .#####
        "00000000", --
        -- 4 
        "00011100", -- ...###
        "00111100", -- ..####
        "01101100", -- .## ##
        "11001100", -- ## .##
        "11111110", -- #######
        "00001100", -- ....##
        "00001100", -- ....##
        "00000000", --
        -- 5 
        "11111100", -- ######
        "11000000", -- ##
        "11111100", -- ######
        "00000110", -- ##
        "00000110", -- ##
        "11000110", -- ## ##
        "01111100", -- #####
        "00000000", --
        -- 6 
        "00111100", -- ####
        "01100000", -- ##
        "11000000", -- ##
        "11111100", -- ######
        "11000110", -- ## ##
        "11000110", -- ## ##
        "01111100", -- #####
        "00000000", --
        -- 7 
        "11111110", -- #######
        "11000110", -- ## ##
        "00001100", -- ##
        "00011000", -- ##
        "00110000", -- ##
        "00110000", -- ##
        "00110000", -- ##
        "00000000", --
        -- 8 
        "01111000", -- .####
        "11000100", -- ## ..#
        "11100100", -- ### .#
        "01111000", -- .####
        "10011110", -- # ####
        "10000110", -- # ..##
        "01111100", -- .#####
        "00000000", --
        -- 9 
        "01111100", -- .#####
        "11000110", -- ##. .##
        "11000110", -- ##. .##
        "01111110", -- .######
        "00000110", -- .....##
        "00001100", -- ....##
        "01111000", -- ####
        "00000000", --
		  -- 10
		  "01111100", -- .#####
        "11111110", -- #######
        "11000110", -- ##...##
        "00001100", -- ....##
        "00111000", -- ..###
        "00000000", --
        "00111000", -- ..###
        "00000000", --
		  -- 11 A
		  "00111000", -- ..###
        "01101100", -- .## ##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11111110", -- #######
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "00000000", --
        -- 12 B
        "11111100", -- ######
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11111100", -- ######
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11111100", -- ######
        "00000000", --
        -- 13
        "00111100", -- ..####
        "01100110", -- .## .##
        "11000000", -- ##
        "11000000", -- ##
        "11000000", -- ##
        "01100110", -- .## .##
        "00111100", -- ..####
        "00000000", --
        -- 14
        "11111000", -- #####
        "11001100", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11001100", -- ## ##
        "11111000", -- #####
        "00000000", --
        -- 15
        "11111110", -- #######
        "11000000", -- ##
        "11000000", -- ##
        "11111100", -- ######
        "11000000", -- ##
        "11000000", -- ##
        "11111110", -- #######
        "00000000", --
        -- 16
        "11111110", -- #######
        "11000000", -- ##
        "11000000", -- ##
        "11111100", -- ######
        "11000000", -- ##
        "11000000", -- ##
        "11000000", -- ##
        "00000000", --
        -- 17
        "00111110", -- #####
        "01100000", -- ##
        "11000000", -- ##
        "11001110", -- ## ###
        "11000110", -- ## ##
        "01100110", -- ## ##
        "00111110", -- #####
        "00000000", --
        -- 13
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11111110", -- #######
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "00000000", --
        -- 24
        "01111110", --. ######
        "00011000", -- ...##
        "00011000", -- ...##
        "00011000", -- ...##
        "00011000", -- ...##
        "00011000", -- ...##
        "01111110", --. ######
        "00000000", --
        -- 25
        "00011110", -- ####
        "00001100", -- ##
        "00001100", -- ##
        "00001100", -- ##
        "00001100", -- ##
        "10001100", -- # ##
        "01111000", -- ####
        "00000000", --
        -- 26
        "11000110", -- ## ##
        "11001100", -- ## ##
        "11011000", -- ## ##
        "11110000", -- ####
        "11111000", -- #####
        "11011100", -- ## ###
        "11001110", -- ## ###
        "00000000", --
        -- 27
        "01100000", -- ##
        "01100000", -- ##
        "01100000", -- ##
        "01100000", -- ##
        "01100000", -- ##
        "01100000", -- ##
        "01111110", -- ######
        "00000000", --
        -- 28
        "11000110", -- ## ##
        "11101110", -- ### ###
        "11111110", -- #######
        "11111110", -- #######
        "11010110", -- ## # ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "00000000", --
        -- 29
        "11000110", -- ## ##
        "11100110", -- ### ##
        "11110110", -- #### ##
        "11111110", -- #######
        "11011110", -- ## ####
        "11001110", -- ## ###
        "11000110", -- ## ##
        "00000000", --
        -- 30
        "01111100", -- .#####
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "11000110", -- ## ..##
        "01111100", -- .#####
        "00000000", --
        -- 31
        "11111100", -- ######
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11111100", -- ######
        "11000000", -- ##
        "11000000", -- ##
        "00000000", --
        -- 32
        "01111100", -- #####
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11011110", -- ## ####
        "11001100", -- ## ##
        "01111010", -- #### #
        "00000000", --
        -- 33
        "11111100", -- ######
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11001110", -- ## ###
        "11111000", -- #####
        "11011100", -- ## ###
        "11001110", -- ## ###
        "00000000", --
        -- 34
        "01111000", -- ####
        "11001100", -- ## ##
        "11000000", -- ##
        "01111100", -- #####
        "00000110", -- ##
        "11000110", -- ## ##
        "01111100", -- #####
        "00000000", --
        -- 35
        "01111110", -- ######
        "00011000", -- ##
        "00011000", -- ##
        "00011000", -- ##
        "00011000", -- ##
        "00011000", -- ##
        "00011000", -- ##
        "00000000", --
        -- 36
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "01111100", -- #####
        "00000000", --
        -- 37
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11101110", -- ### ###
        "01111100", -- #####
        "00111000", -- ###
        "00010000", -- #
        "00000000", --
        -- 38
        "11000110", -- ## ##
        "11000110", -- ## ##
        "11010110", -- ## # ##
        "11111110", -- #######
        "11111110", -- #######
        "11101110", -- ### ###
        "11000110", -- ## ##
        "00000000", --
        -- 39
        "11000110", -- ##...##
        "11101110", -- ### ###
        "01111100", -- .#####
        "00111000", -- ..###
        "01111100", -- .#####
        "11101110", -- ### ###
        "11000110", -- ##...##
        "00000000", --
        -- 40
        "01100110", -- ## ##
        "01100110", -- ## ##
        "01100110", -- ## ##
        "00111100", -- ####
        "00011000", -- ##
        "00011000", -- ##
        "00011000", -- ##
        "00000000", --
        -- 41
        "11111110", -- #######
        "00001110", -- ....##
        "00011100", -- ...###
        "00111000", -- ..###
        "01110000", -- .###
        "11100000", -- ###
        "11111110", -- #######
        "00000000", --
         -- 42
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        -- 43
        "00111000", -- ###
        "00111000", -- ###
        "00111000", -- ###
        "00110000", -- ##
        "00110000", -- ##
        "00000000", --
        "00110000", -- ##
        "00000000", --
        -- 44
        "00000000", --
        "00000000", --
        "00000000", --
        "01111100", -- #####
        "00000000", --
        "00000000", --
        "00000000", --
        "00000000", --
        -- 45
        "00000000", --
        "00110000", -- ##
        "00110000", -- ##
        "00000000", -- 
        "00000000", --
        "00110000", -- ##
        "00110000", -- ##
        "00000000", --
        -- 46
        "00100000", -- #
        "00110000", -- ##
        "00111000", -- ###
        "00111100", -- ####
        "00111000", -- ###
        "00110000", -- ##
        "00100000", -- #
        "00000000" --
    );
begin
    data <= FONT(conv_integer(addr));
end content;